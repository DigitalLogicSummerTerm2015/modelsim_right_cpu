`timescale 1ns/1ps

module ROM(addr, data);
input [31:0] addr;
output [31:0] data;

localparam ROM_SIZE = 32;

reg [31:0] data;
reg [31:0] ROM_DATA[ROM_SIZE-1:0];

always@(*)
    case(addr[9:2])  // Address Must Be Word Aligned.
        0: data <= 32'h08000003;
        1: data <= 32'h08000032;
        2: data <= 32'h08000070;
        3: data <= 32'h200800c0;
        4: data <= 32'hac080000;
        5: data <= 32'h200800f9;
        6: data <= 32'hac080004;
        7: data <= 32'h200800a4;
        8: data <= 32'hac080008;
        9: data <= 32'h200800b0;
        10: data <= 32'hac08000c;
        11: data <= 32'h20080099;
        12: data <= 32'hac080010;
        13: data <= 32'h20080092;
        14: data <= 32'hac080014;
        15: data <= 32'h20080082;
        16: data <= 32'hac080018;
        17: data <= 32'h200800f8;
        18: data <= 32'hac08001c;
        19: data <= 32'h20080080;
        20: data <= 32'hac080020;
        21: data <= 32'h20080090;
        22: data <= 32'hac080024;
        23: data <= 32'h20080088;
        24: data <= 32'hac080028;
        25: data <= 32'h20080083;
        26: data <= 32'hac08002c;
        27: data <= 32'h200800c6;
        28: data <= 32'hac080030;
        29: data <= 32'h200800a1;
        30: data <= 32'hac080034;
        31: data <= 32'h20080086;
        32: data <= 32'hac080038;
        33: data <= 32'h2008008e;
        34: data <= 32'hac08003c;
        35: data <= 32'h3c174000;
        36: data <= 32'haee00008;
        37: data <= 32'h20088000;
        38: data <= 32'haee80000;
        39: data <= 32'h2008ffff;
        40: data <= 32'haee80004;
        41: data <= 32'h0c00002a;
        42: data <= 32'h3c088000;
        43: data <= 32'h01004027;
        44: data <= 32'h011ff824;
        45: data <= 32'h23ff0014;
        46: data <= 32'h03e00008;
        47: data <= 32'h20080003;
        48: data <= 32'haee80008;
        49: data <= 32'h08000031;
        50: data <= 32'h3c174000;
        51: data <= 32'h8ee80008;
        52: data <= 32'h2009fff9;
        53: data <= 32'h01094024;
        54: data <= 32'haee80008;
        55: data <= 32'h8ee80020;
        56: data <= 32'h11000018;
        57: data <= 32'h8ee40018;
        58: data <= 32'h8ee5001c;
        59: data <= 32'h1080000d;
        60: data <= 32'h10a0000e;
        61: data <= 32'h00808020;
        62: data <= 32'h00a08820;
        63: data <= 32'h0211402a;
        64: data <= 32'h15000002;
        65: data <= 32'h02118022;
        66: data <= 32'h0800003f;
        67: data <= 32'h02004020;
        68: data <= 32'h02208020;
        69: data <= 32'h01008820;
        70: data <= 32'h1620fff8;
        71: data <= 32'h02001020;
        72: data <= 32'h0800004c;
        73: data <= 32'h00051020;
        74: data <= 32'h0800004c;
        75: data <= 32'h00041020;
        76: data <= 32'haee20024;
        77: data <= 32'h20080001;
        78: data <= 32'haee80028;
        79: data <= 32'haee00028;
        80: data <= 32'haee2000c;
        81: data <= 32'h8eec0014;
        82: data <= 32'h000c6202;
        83: data <= 32'h000c6040;
        84: data <= 32'h218c0001;
        85: data <= 32'h318c000f;
        86: data <= 32'h2009000d;
        87: data <= 32'h200a000b;
        88: data <= 32'h200b0007;
        89: data <= 32'h11890005;
        90: data <= 32'h118a0006;
        91: data <= 32'h118b0007;
        92: data <= 32'h200c000e;
        93: data <= 32'h00a06820;
        94: data <= 32'h08000065;
        95: data <= 32'h00056902;
        96: data <= 32'h08000065;
        97: data <= 32'h00806820;
        98: data <= 32'h08000065;
        99: data <= 32'h00046902;
        100: data <= 32'h08000065;
        101: data <= 32'h31ad000f;
        102: data <= 32'h000d6880;
        103: data <= 32'h8dad0000;
        104: data <= 32'h000c6200;
        105: data <= 32'h018d4020;
        106: data <= 32'haee80014;
        107: data <= 32'h8ee80008;
        108: data <= 32'h20090002;
        109: data <= 32'h01094025;
        110: data <= 32'haee80008;
        111: data <= 32'h03400008;
        112: data <= 32'h03400008;
        default: data <= 32'h0800_0000;
    endcase
endmodule

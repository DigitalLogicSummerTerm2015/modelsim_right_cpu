`timescale 1ns/1ps

module ROM(addr, data);
input [31:0] addr;
output [31:0] data;

localparam ROM_SIZE = 32;

reg [31:0] data;
reg [31:0] ROM_DATA[ROM_SIZE-1:0];

always@(*)
    case(addr[9:2])  // Address Must Be Word Aligned.
        0: data <= 32'h08000003;
        1: data <= 32'h08000032;
        2: data <= 32'h08000087;
        3: data <= 32'h20080040;
        4: data <= 32'hac080000;
        5: data <= 32'h20080079;
        6: data <= 32'hac080004;
        7: data <= 32'h20080024;
        8: data <= 32'hac080008;
        9: data <= 32'h20080030;
        10: data <= 32'hac08000c;
        11: data <= 32'h20080019;
        12: data <= 32'hac080010;
        13: data <= 32'h20080012;
        14: data <= 32'hac080014;
        15: data <= 32'h20080002;
        16: data <= 32'hac080018;
        17: data <= 32'h20080078;
        18: data <= 32'hac08001c;
        19: data <= 32'h20080000;
        20: data <= 32'hac080020;
        21: data <= 32'h20080010;
        22: data <= 32'hac080024;
        23: data <= 32'h20080008;
        24: data <= 32'hac080028;
        25: data <= 32'h20080003;
        26: data <= 32'hac08002c;
        27: data <= 32'h20080046;
        28: data <= 32'hac080030;
        29: data <= 32'h20080021;
        30: data <= 32'hac080034;
        31: data <= 32'h20080006;
        32: data <= 32'hac080038;
        33: data <= 32'h2008000e;
        34: data <= 32'hac08003c;
        35: data <= 32'h3c174000;
        36: data <= 32'haee00008;
        37: data <= 32'h20088000;
        38: data <= 32'haee80000;
        39: data <= 32'h2008ffff;
        40: data <= 32'haee80004;
        41: data <= 32'h0c00002a;
        42: data <= 32'h3c088000;
        43: data <= 32'h01004027;
        44: data <= 32'h011ff824;
        45: data <= 32'h23ff0014;
        46: data <= 32'h03e00008;
        47: data <= 32'h20080003;
        48: data <= 32'haee80008;
        49: data <= 32'h08000031;
        50: data <= 32'h3c174000;
        51: data <= 32'h8ee80008;
        52: data <= 32'h2009fff9;
        53: data <= 32'h01094024;
        54: data <= 32'h00000000;
        55: data <= 32'h00000000;
        56: data <= 32'h00000000;
        57: data <= 32'haee80008;
        58: data <= 32'h00000000;
        59: data <= 32'h00000000;
        60: data <= 32'h00000000;
        61: data <= 32'h8ee80020;
        62: data <= 32'h00000000;
        63: data <= 32'h00000000;
        64: data <= 32'h00000000;
        65: data <= 32'h11000024;
        66: data <= 32'h00000000;
        67: data <= 32'h00000000;
        68: data <= 32'h00000000;
        69: data <= 32'h8ee40018;
        70: data <= 32'h00000000;
        71: data <= 32'h00000000;
        72: data <= 32'h00000000;
        73: data <= 32'h8ee5001c;
        74: data <= 32'h00000000;
        75: data <= 32'h00000000;
        76: data <= 32'h00000000;
        77: data <= 32'h10800017;
        78: data <= 32'h00000000;
        79: data <= 32'h00000000;
        80: data <= 32'h00000000;
        81: data <= 32'h10a00013;
        82: data <= 32'h00000000;
        83: data <= 32'h00000000;
        84: data <= 32'h00000000;
        85: data <= 32'h00808020;
        86: data <= 32'h00a08820;
        87: data <= 32'h0211402a;
        88: data <= 32'h15000002;
        89: data <= 32'h02118022;
        90: data <= 32'h08000057;
        91: data <= 32'h02004020;
        92: data <= 32'h02208020;
        93: data <= 32'h01008820;
        94: data <= 32'h1620fff8;
        95: data <= 32'h02001020;
        96: data <= 32'haee20024;
        97: data <= 32'h20080001;
        98: data <= 32'haee80028;
        99: data <= 32'haee00028;
        100: data <= 32'h08000066;
        101: data <= 32'h00001020;
        102: data <= 32'haee2000c;
        103: data <= 32'h8eec0014;
        104: data <= 32'h000c6202;
        105: data <= 32'h318c000f;
        106: data <= 32'h000c6040;
        107: data <= 32'h20080001;
        108: data <= 32'h20090002;
        109: data <= 32'h200a0004;
        110: data <= 32'h200b0008;
        111: data <= 32'h11880004;
        112: data <= 32'h11890005;
        113: data <= 32'h118a0006;
        114: data <= 32'h118b0007;
        115: data <= 32'h200c0001;
        116: data <= 32'h00046902;
        117: data <= 32'h0800007c;
        118: data <= 32'h00806820;
        119: data <= 32'h0800007c;
        120: data <= 32'h00056902;
        121: data <= 32'h0800007c;
        122: data <= 32'h00a06820;
        123: data <= 32'h0800007c;
        124: data <= 32'h31ad000f;
        125: data <= 32'h000d6880;
        126: data <= 32'h8dad0000;
        127: data <= 32'h000c6200;
        128: data <= 32'h018d4020;
        129: data <= 32'haee80014;
        130: data <= 32'h8ee80008;
        131: data <= 32'h20090002;
        132: data <= 32'h01094025;
        133: data <= 32'haee80008;
        134: data <= 32'h03400008;
        135: data <= 32'h03400008;
        default: data <= 32'h0800_0000;
    endcase
endmodule

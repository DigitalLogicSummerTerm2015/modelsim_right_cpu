`timescale 1ns/1ps

module ROM(addr, data);
input [31:0] addr;
output [31:0] data;

localparam ROM_SIZE = 32;

reg [31:0] data;
reg [31:0] ROM_DATA[ROM_SIZE-1:0];

always@(*)
    case(addr[9:2])  // Address Must Be Word Aligned.
        0: data <= 32'h08000003;
        1: data <= 32'h08000044;
        2: data <= 32'h080000be;
        3: data <= 32'h200800c0;
        4: data <= 32'hac080000;
        5: data <= 32'h200800f9;
        6: data <= 32'hac080004;
        7: data <= 32'h200800a4;
        8: data <= 32'hac080008;
        9: data <= 32'h200800b0;
        10: data <= 32'hac08000c;
        11: data <= 32'h20080099;
        12: data <= 32'hac080010;
        13: data <= 32'h20080092;
        14: data <= 32'hac080014;
        15: data <= 32'h20080082;
        16: data <= 32'hac080018;
        17: data <= 32'h200800f8;
        18: data <= 32'hac08001c;
        19: data <= 32'h20080080;
        20: data <= 32'hac080020;
        21: data <= 32'h20080090;
        22: data <= 32'hac080024;
        23: data <= 32'h20080088;
        24: data <= 32'hac080028;
        25: data <= 32'h20080083;
        26: data <= 32'hac08002c;
        27: data <= 32'h200800c6;
        28: data <= 32'hac080030;
        29: data <= 32'h200800a1;
        30: data <= 32'hac080034;
        31: data <= 32'h20080086;
        32: data <= 32'hac080038;
        33: data <= 32'h2008008e;
        34: data <= 32'hac08003c;
        35: data <= 32'h3c174000;
        36: data <= 32'haee00008;
        37: data <= 32'h20088000;
        38: data <= 32'h00000000;
        39: data <= 32'h00000000;
        40: data <= 32'h00000000;
        41: data <= 32'haee80000;
        42: data <= 32'h00000000;
        43: data <= 32'h00000000;
        44: data <= 32'h00000000;
        45: data <= 32'h2008ffff;
        46: data <= 32'h00000000;
        47: data <= 32'h00000000;
        48: data <= 32'h00000000;
        49: data <= 32'haee80004;
        50: data <= 32'h00000000;
        51: data <= 32'h00000000;
        52: data <= 32'h00000000;
        53: data <= 32'h0c000036;
        54: data <= 32'h3c088000;
        55: data <= 32'h01004027;
        56: data <= 32'h011ff824;
        57: data <= 32'h23ff0014;
        58: data <= 32'h03e00008;
        59: data <= 32'h20080003;
        60: data <= 32'h00000000;
        61: data <= 32'h00000000;
        62: data <= 32'h00000000;
        63: data <= 32'haee80008;
        64: data <= 32'h00000000;
        65: data <= 32'h00000000;
        66: data <= 32'h00000000;
        67: data <= 32'h08000043;
        68: data <= 32'h3c174000;
        69: data <= 32'h00000000;
        70: data <= 32'h00000000;
        71: data <= 32'h00000000;
        72: data <= 32'h8ee80008;
        73: data <= 32'h00000000;
        74: data <= 32'h00000000;
        75: data <= 32'h00000000;
        76: data <= 32'h2009fff9;
        77: data <= 32'h01094024;
        78: data <= 32'h00000000;
        79: data <= 32'h00000000;
        80: data <= 32'h00000000;
        81: data <= 32'haee80008;
        82: data <= 32'h00000000;
        83: data <= 32'h00000000;
        84: data <= 32'h00000000;
        85: data <= 32'h8ee80020;
        86: data <= 32'h00000000;
        87: data <= 32'h00000000;
        88: data <= 32'h00000000;
        89: data <= 32'h1100002d;
        90: data <= 32'h00000000;
        91: data <= 32'h00000000;
        92: data <= 32'h00000000;
        93: data <= 32'h8ee40018;
        94: data <= 32'h00000000;
        95: data <= 32'h00000000;
        96: data <= 32'h00000000;
        97: data <= 32'h8ee5001c;
        98: data <= 32'h00000000;
        99: data <= 32'h00000000;
        100: data <= 32'h00000000;
        101: data <= 32'h1080000d;
        102: data <= 32'h10a0000e;
        103: data <= 32'h00808020;
        104: data <= 32'h00a08820;
        105: data <= 32'h0211402a;
        106: data <= 32'h15000002;
        107: data <= 32'h02118022;
        108: data <= 32'h08000069;
        109: data <= 32'h02004020;
        110: data <= 32'h02208020;
        111: data <= 32'h01008820;
        112: data <= 32'h1620fff8;
        113: data <= 32'h02001020;
        114: data <= 32'h08000076;
        115: data <= 32'h00051020;
        116: data <= 32'h08000076;
        117: data <= 32'h00041020;
        118: data <= 32'h00000000;
        119: data <= 32'h00000000;
        120: data <= 32'h00000000;
        121: data <= 32'haee20024;
        122: data <= 32'h20080001;
        123: data <= 32'h00000000;
        124: data <= 32'h00000000;
        125: data <= 32'h00000000;
        126: data <= 32'haee80028;
        127: data <= 32'h00000000;
        128: data <= 32'h00000000;
        129: data <= 32'h00000000;
        130: data <= 32'haee00028;
        131: data <= 32'h00000000;
        132: data <= 32'h00000000;
        133: data <= 32'h00000000;
        134: data <= 32'haee2000c;
        135: data <= 32'h00000000;
        136: data <= 32'h00000000;
        137: data <= 32'h00000000;
        138: data <= 32'h8eec0014;
        139: data <= 32'h00000000;
        140: data <= 32'h00000000;
        141: data <= 32'h00000000;
        142: data <= 32'h000c6202;
        143: data <= 32'h000c6040;
        144: data <= 32'h218c0001;
        145: data <= 32'h318c000f;
        146: data <= 32'h2009000d;
        147: data <= 32'h200a000b;
        148: data <= 32'h200b0007;
        149: data <= 32'h11890005;
        150: data <= 32'h118a0006;
        151: data <= 32'h118b0007;
        152: data <= 32'h200c000e;
        153: data <= 32'h00a06820;
        154: data <= 32'h080000a1;
        155: data <= 32'h00056902;
        156: data <= 32'h080000a1;
        157: data <= 32'h00806820;
        158: data <= 32'h080000a1;
        159: data <= 32'h00046902;
        160: data <= 32'h080000a1;
        161: data <= 32'h31ad000f;
        162: data <= 32'h000d6880;
        163: data <= 32'h8dad0000;
        164: data <= 32'h00000000;
        165: data <= 32'h00000000;
        166: data <= 32'h00000000;
        167: data <= 32'h000c6200;
        168: data <= 32'h018d4020;
        169: data <= 32'h00000000;
        170: data <= 32'h00000000;
        171: data <= 32'h00000000;
        172: data <= 32'haee80014;
        173: data <= 32'h00000000;
        174: data <= 32'h00000000;
        175: data <= 32'h00000000;
        176: data <= 32'h8ee80008;
        177: data <= 32'h00000000;
        178: data <= 32'h00000000;
        179: data <= 32'h00000000;
        180: data <= 32'h20090002;
        181: data <= 32'h01094025;
        182: data <= 32'h00000000;
        183: data <= 32'h00000000;
        184: data <= 32'h00000000;
        185: data <= 32'haee80008;
        186: data <= 32'h00000000;
        187: data <= 32'h00000000;
        188: data <= 32'h00000000;
        189: data <= 32'h03400008;
        190: data <= 32'h03400008;
        default: data <= 32'h0800_0000;
    endcase
endmodule
